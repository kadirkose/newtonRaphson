library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;	
use ieee.std_logic_unsigned.all;	

entity newton_raphson is
	generic(	
		DATA_WIDTH 				: in 	natural := 32;												 	-- RAM dimensions
		ADDR_WIDTH 				: in 	natural := 128;								
		CLK_FREQ      			: in 	integer := 125e6;   											-- set system clock frequency in Hz
		BAUD_RATE     			: in 	integer := 115200;   										-- baud rate value
		PARITY_BIT    			: in 	string  := "none"; 											-- legal values: "none", "even", "odd", "mark", "space"
		USE_DEBOUNCER 			: in 	boolean := false   											-- enable/disable debouncer		
	);
	port(
		clk						: in 		std_logic;
		reset						: in 		std_logic;
		UART_TXD   				: out 	std_logic;
		UART_RXD   				: in  	std_logic;
		leds						: out 	std_logic_vector(9 downto 0):= (others => '0');	-- these connected to terasIC DE10-Lite LED pins
		ledg						: out 	std_logic_vector(7 downto 0):= (others => '0')
	);
end newton_raphson;

architecture logic of newton_raphson is
	
	component calculator_rtl
		port(
			ledg								: out std_logic_vector(7 downto 0):= (others => '0');
			clk								: in 	std_logic;
			reset								: in 	std_logic;
			start_op							: in 	std_logic;
			degree							: in 	integer;
			degree_min						: in 	integer;
			variable_value					: in	std_logic_vector(31 downto 0):= (others => '0');
			op_result						: out	std_logic_vector(31 downto 0):= (others => '0');
			complete_op_flag				: out	std_logic:= '0';
			error_value						: out std_logic_vector(31 downto 0):= (others => '0');
			float_in0        				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in1        				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in2        				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in3        				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in4        				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in5        				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in6        				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in7        				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in8        				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in9        				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in10						: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in11       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in12       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in13       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in14       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in15       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in16       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in17       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in18       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in19       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in20       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in21       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in22       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in23       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in24       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in25       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in26       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in27       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in28       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in29       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in30       				: in 	std_logic_vector(31 downto 0):= (others => '0');
			float_in31       				: in 	std_logic_vector(31 downto 0):= (others => '0')
		);
	end component;
	
	component uart
		generic(
			CLK_FREQ      				: in 	integer := 125e6;   									-- system clock frequency in Hz
			BAUD_RATE     				: in 	integer := 115200; 									-- baud rate value
			PARITY_BIT    				: in 	string  := "none"; 									-- type of parity: "none", "even", "odd", "mark", "space"
			USE_DEBOUNCER 				: in 	boolean := FALSE   									-- enable/disable debouncer
		);
		port(
			-- CLOCK AND RESET
			CLK         				: in  std_logic; 												-- system clock
			RST         				: in  std_logic; 												-- high active synchronous reset
			-- UART INTERFACE
			UART_TXD    				: out std_logic; 												-- serial transmit data
			UART_RXD    				: in  std_logic; 												-- serial receive data
			-- USER DATA INPUT INTERFACE
			DIN         				: in  std_logic_vector(7 downto 0); 					-- input data to be transmitted over UART
			DIN_VLD     				: in  std_logic; 												-- when DIN_VLD = 1, input data (DIN) are valid
			DIN_RDY     				: out std_logic; 												-- when DIN_RDY = 1, transmitter is ready and valid input data will be accepted for transmiting
			-- USER DATA OUTPUT INTERFACE
			DOUT        				: out std_logic_vector(7 downto 0); 					-- output data received via UART
			DOUT_VLD    				: out std_logic; 												-- when v = 1, output data (DOUT) are valid (is assert only for one clock cycle)
			FRAME_ERROR 				: out std_logic;  											-- when FRAME_ERROR = 1, stop bit was invalid (is assert only for one clock cycle)
			PARITY_ERROR 				: out std_logic  												-- when PARITY_ERROR = 1, parity bit was invalid (is assert only for one clock cycl
		);
	end component;
	
	component fp_comparator
		port (
			a 						: in std_logic_vector(31 downto 0);  -- float32_m23
			b 						: in std_logic_vector(31 downto 0);  -- float32_m23
			q 						: out std_logic_vector(0 downto 0);  -- ufix1
			clk 					: in std_logic;
			areset 				: in std_logic
		);
	end component;
	
	component ip_core_operation_wait is
		port(
			clk					: in 	std_logic;
			ip_wait_reset		: in 	std_logic;
			ip_op_wait_ok		: out std_logic;
			ip_op_wait			: in	std_logic_vector(2 downto 0):= "000"
		);
	end component;

	signal cnt									: integer range 0 to 100:= 0;
	signal count								: integer:= 0;
	signal cycle_count						: std_logic_vector(31 downto 0):= (others => '0');
	signal total_cycle_count				: std_logic_vector(31 downto 0):= (others => '0');

	
	signal u_data_in, u_data_out			: std_logic_vector(7 downto 0);					-- internal UART signals 
	signal u_valid_out, u_valid_in		: std_logic:='0';
	signal u_data_in_ready 					: std_logic:='1';
	signal u_data_in_ready_prev			: std_logic:='1';
	
	signal variable_value					: std_logic_vector(31 downto 0):= (others => '0');

	signal degree_min, degree_max, degree	: integer:= 0;
	
	signal start_opr							: std_logic:= '0';
	signal complete_calculator_flag		: std_logic:= '0';
	signal calculator_result				: std_logic_vector(31 downto 0);
	signal newton_raphson_result			: std_logic_vector(31 downto 0); 
	
	type float32 is array(31 downto 0) of std_logic_vector(31 downto 0);
	signal float_in		: float32:= (others => "00000000000000000000000000000000");
	
	signal float_comp_in1			: std_logic_vector(31 downto 0):= (others => '0');
	signal error_value				: std_logic_vector(31 downto 0):= (others => '0');
	signal float_comp_out			: std_logic_vector(0 downto 0) := (others => '0');
	signal iteration_count			: std_logic_vector(31 downto 0):= (others => '0');
	signal error_const_value		: std_logic_vector(31 downto 0):= (others => '0');
	signal float_comp_in2			: std_logic_vector(31 downto 0):= (others => '0');
	signal interation_limit			: std_logic_vector(31 downto 0):= (others => '0');
	
	signal ip_wait_reset				: std_logic;
	signal ip_op_wait_ok				: std_logic;
	signal ip_op_wait					: std_logic_vector(2 downto 0):= "000";

	
	type machine is(
		get_min_degree, 
		get_max_degree,
		degree_range_control,
		get_var_val, 
		get_error_val,
		get_iteration_val,
		get_coefficients, 
		initialize_calculator,
		complete_calculator, 
		initialize_compare,
		wait_compare,
		complete_compare,
		send_result,
		power_off,
		reset_all_variable,
		idle
	);
	signal state: machine:= get_min_degree;																-- state machine instruction
	
	begin
	
	calculator_block: calculator_rtl
	port map(
	ledg => ledg,
		clk								=> clk,
		reset								=> reset,
		start_op							=> start_opr,
		degree							=> degree,
		degree_min						=> degree_min,
		variable_value					=> variable_value,
		op_result						=> calculator_result,
		error_value						=> error_value,
		complete_op_flag				=> complete_calculator_flag,
		float_in0        				=> float_in(0),  
		float_in1        				=> float_in(1),    
		float_in2        				=> float_in(2),    
		float_in3        				=> float_in(3),    
		float_in4        				=> float_in(4),    
		float_in5        				=> float_in(5),     
		float_in6        				=> float_in(6),    
		float_in7        				=> float_in(7),    
		float_in8        				=> float_in(8),    
		float_in9        				=> float_in(9),    
		float_in10						=> float_in(10),	
		float_in11       				=> float_in(11),   
		float_in12       				=> float_in(12),   
		float_in13       				=> float_in(13),   
		float_in14       				=> float_in(14),   
		float_in15       				=> float_in(15),   
		float_in16       				=> float_in(16),   
		float_in17       				=> float_in(17),   
		float_in18       				=> float_in(18),   
		float_in19       				=> float_in(19),   
		float_in20       				=> float_in(20),   
		float_in21       				=> float_in(21),   
		float_in22       				=> float_in(22),   
		float_in23       				=> float_in(23),   
		float_in24       				=> float_in(24),   
		float_in25       				=> float_in(25),   
		float_in26       				=> float_in(26),   
		float_in27       				=> float_in(27),   
		float_in28       				=> float_in(28),   
		float_in29       				=> float_in(29),   
		float_in30       				=> float_in(30),   
		float_in31       				=> float_in(31)
	);
	
	uart_block: uart
   generic map(
       CLK_FREQ      => CLK_FREQ,
       BAUD_RATE     => BAUD_RATE,
       PARITY_BIT    => PARITY_BIT,
       USE_DEBOUNCER => USE_DEBOUNCER
   )
   port map(
       CLK         	=> clk,
       RST         	=> not reset,																	-- UART module reset is reverse
       -- UART INTERFACE
       UART_TXD    	=> UART_TXD,
       UART_RXD    	=> UART_RXD,
       -- USER DATA OUTPUT INTERFACE
       DOUT        	=> u_data_out,
       DOUT_VLD    	=> u_valid_out,
       FRAME_ERROR 	=> open,
		 PARITY_ERROR	=> open,
       -- USER DATA INPUT INTERFACE
       DIN         	=> u_data_in,
       DIN_VLD     	=> u_valid_in,
       DIN_RDY     	=> u_data_in_ready
   );
	
	float_comparator_block: fp_comparator
	port map(
		clk    => clk,
		areset => not reset,
		a      => float_comp_in1,
		b      => float_comp_in2,
		q      => float_comp_out
	);
	
	ip_core_wait_block: ip_core_operation_wait
	port map(
		clk				=> clk,
		ip_wait_reset	=> ip_wait_reset,
		ip_op_wait_ok	=> ip_op_wait_ok,
		ip_op_wait		=> ip_op_wait
	);		
	
	process(clk, reset)
	begin
		if(reset = '0') then
			u_valid_in 					<= '0';
			u_data_in 					<= "01010010";														-- ASCII 'R'
			cnt 							<= 0;
			count							<= 0;
			cycle_count					<= (others => '0');
			total_cycle_count			<= (others => '0');
			state 						<= idle;
			degree_min					<= 0;	
			degree_max					<= 0;	
			degree						<= 0;	
			start_opr					<= '0';			
			leds 							<= "0000000000";
			variable_value		  		<= (others => '0');
			float_in(0)  				<= (others => '0');
			float_in(1)  				<= (others => '0');
			float_in(2)  				<= (others => '0');
			float_in(3)  				<= (others => '0');
			float_in(4)  				<= (others => '0');
			float_in(5)  				<= (others => '0');
			float_in(6) 				<= (others => '0');
			float_in(7)  				<= (others => '0');
			float_in(8)  				<= (others => '0');
			float_in(9)  				<= (others => '0');
			float_in(10)  				<= (others => '0');
			float_in(11)				<= (others => '0');
			float_in(12)  				<= (others => '0');
			float_in(13)  				<= (others => '0');
			float_in(14)  				<= (others => '0');
			float_in(15)  				<= (others => '0');
			float_in(16)  				<= (others => '0');
			float_in(17)  				<= (others => '0');
			float_in(18) 				<= (others => '0');
			float_in(19)  				<= (others => '0');
			float_in(20)  				<= (others => '0');
			float_in(21)  				<= (others => '0');
			float_in(22)  				<= (others => '0');
			float_in(23)  				<= (others => '0');
			float_in(24)  				<= (others => '0');
			float_in(25)  				<= (others => '0');
			float_in(26)  				<= (others => '0');
			float_in(27)  				<= (others => '0');
			float_in(28)  				<= (others => '0');
			float_in(29)  				<= (others => '0');
			float_in(30)  				<= (others => '0');
			float_in(31)  				<= (others => '0');
			iteration_count			<= (others => '0');
			error_const_value			<= (others => '0');
			interation_limit			<= (others => '0');
			float_comp_in1				<= (others => '0');
		elsif(rising_edge(clk)) then
			u_data_in_ready_prev <= u_data_in_ready;
			case state is
			
				when idle =>
					leds	 		<= "1111111111";
					u_valid_in 					<= '0';
					u_data_in 					<= "01010010";														-- ASCII 'R'
					cnt 							<= 0;
					count							<= 0;
					cycle_count					<= (others => '0');
					total_cycle_count			<= (others => '0');
					state 						<= idle;
					degree_min					<= 0;	
					degree_max					<= 0;	
					degree						<= 0;	
					start_opr					<= '0';			
					variable_value		  		<= (others => '0');
					float_in(0)  				<= (others => '0');
					float_in(1)  				<= (others => '0');
					float_in(2)  				<= (others => '0');
					float_in(3)  				<= (others => '0');
					float_in(4)  				<= (others => '0');
					float_in(5)  				<= (others => '0');
					float_in(6) 				<= (others => '0');
					float_in(7)  				<= (others => '0');
					float_in(8)  				<= (others => '0');
					float_in(9)  				<= (others => '0');
					float_in(10)  				<= (others => '0');
					float_in(11)				<= (others => '0');
					float_in(12)  				<= (others => '0');
					float_in(13)  				<= (others => '0');
					float_in(14)  				<= (others => '0');
					float_in(15)  				<= (others => '0');
					float_in(16)  				<= (others => '0');
					float_in(17)  				<= (others => '0');
					float_in(18) 				<= (others => '0');
					float_in(19)  				<= (others => '0');
					float_in(20)  				<= (others => '0');
					float_in(21)  				<= (others => '0');
					float_in(22)  				<= (others => '0');
					float_in(23)  				<= (others => '0');
					float_in(24)  				<= (others => '0');
					float_in(25)  				<= (others => '0');
					float_in(26)  				<= (others => '0');
					float_in(27)  				<= (others => '0');
					float_in(28)  				<= (others => '0');
					float_in(29)  				<= (others => '0');
					float_in(30)  				<= (others => '0');
					float_in(31)  				<= (others => '0');
					iteration_count			<= (others => '0');
					error_const_value			<= (others => '0');
					interation_limit			<= (others => '0');
					float_comp_in1				<= (others => '0');
					start_opr	<= '0';
					if(u_valid_out = '1') then																-- if data came from UART
						state 	<= get_min_degree;
					end if;
			
				when get_min_degree =>
					leds	 		<= "0000000001";
					total_cycle_count <= total_cycle_count + 1;
					degree_min 	<= to_integer(unsigned(u_data_out));
					if(to_integer(unsigned(u_data_out)) > 31) then
						state 	<= idle;
					else
						state 	<= get_max_degree;
					end if;
					
				when get_max_degree =>
					total_cycle_count <= total_cycle_count + 1;
					leds	 		<= "0000000010";
					if(u_valid_out = '1') then																-- if data came from UART
						degree_max 	<= to_integer(unsigned(u_data_out));
						if(to_integer(unsigned(u_data_out)) > 31) then
							state 	<= idle;
						else
							state 	<= degree_range_control;
						end if;
					end if;	
					
				when degree_range_control =>
					total_cycle_count <= total_cycle_count + 1;
					leds	 		<= "0000000100";
					if(degree_min + degree_max > 31) then												-- degree must be in range [-31,31] with maximum 32 coefficients
						state 	<= idle;
					else
						state 	<= get_var_val;
						degree 	<= degree_max + degree_min + 1;
					end if;
					
					
				when get_var_val =>
					total_cycle_count <= total_cycle_count + 1;
					leds	 		<= "0000001000";
					if(u_valid_out = '1') then																-- if data came from UART	
						cnt 		<= (cnt + 1);
						variable_value((31 - cnt*8) downto (24 - cnt*8)) <= u_data_out;
						if(cnt = 3) then
							cnt 			<= 0;
							state 		<= get_error_val;
						end if;
					end if;
					
				when get_error_val =>
					total_cycle_count <= total_cycle_count + 1;
					leds	 		<= "0000010000";
					if(u_valid_out = '1') then																-- if data came from UART	
						cnt 		<= (cnt + 1);
						error_const_value((31 - cnt*8) downto (24 - cnt*8)) <= u_data_out;
						if(cnt = 3) then
							cnt 			<= 0;
							state 		<= get_iteration_val;
						end if;
					end if;
					
				when get_iteration_val =>
					total_cycle_count <= total_cycle_count + 1;
					leds	 		<= "0000100000";
					if(u_valid_out = '1') then																-- if data came from UART	
						cnt 		<= (cnt + 1);
						interation_limit((31 - cnt*8) downto (24 - cnt*8)) <= u_data_out;
						if(cnt = 3) then
							cnt 			<= 0;
							state 		<= get_coefficients;
						end if;
					end if;
					
				when get_coefficients =>
					total_cycle_count <= total_cycle_count + 1;
					leds	 		<= "0001000000";
					if(cnt = 4) then
						count 		<= (count + 1);
						cnt 			<= 0;
						if(count = degree - 1) then														-- end of given degree
							state 	<= initialize_calculator;
							count 	<= 0;
						end if;
					end if;
					
					if(u_valid_out = '1') then																-- if data came from UART	
						cnt 			<= (cnt + 1);
						float_in(count)((31 - cnt*8) downto (24 - cnt*8)) <= u_data_out;
					end if;
					
				when initialize_calculator =>
					iteration_count <= iteration_count + 1;
					cycle_count <= cycle_count + 1;
					total_cycle_count <= total_cycle_count + 1;
					leds	 		<= "0010000000";
					start_opr 	<= '1';
					state 		<= complete_calculator;
					
				when complete_calculator =>
					leds	 				<= "0100000000";			
					total_cycle_count <= total_cycle_count + 1;
					cycle_count <= cycle_count + 1;
					if(complete_calculator_flag = '1') then
						state 		<= initialize_compare;
						start_opr 	<= '0';
						newton_raphson_result <= calculator_result;
					end if;
					
				when initialize_compare =>
					float_comp_in1 		<= error_value;
					float_comp_in2			<= error_const_value;
					float_comp_in1(31)	<= '0';
					cycle_count <= cycle_count + 1;
					total_cycle_count <= total_cycle_count + 1;
					leds	 				<= "0100000001";	
					ip_op_wait				<= "101";											-- karşılaştırma bekleme kodu
					ip_wait_reset			<= '1';
					state <= wait_compare;

				when wait_compare =>
					total_cycle_count <= total_cycle_count + 1;
					cycle_count <= cycle_count + 1;
					if(ip_op_wait_ok= '1') then
						ip_op_wait			<= "000";
						ip_wait_reset		<= '0';
						state 				<= complete_compare;
					end if;
					
				when complete_compare =>
					cycle_count <= cycle_count + 1;
					total_cycle_count <= total_cycle_count + 1;
					leds	 				<= "1000000001";	
					if(iteration_count < (interation_limit + 1)) then
						if(float_comp_out = "0" ) then
							state <= initialize_calculator;
							variable_value <= newton_raphson_result;
						else
							state <= send_result;
						end if;
					else
						state <= send_result;
					end if;
					
				when send_result =>
					leds	 		<= "1000000010";
					total_cycle_count <= total_cycle_count + 1;
					u_valid_in 	<= '0';
					if(u_data_in_ready = '0' and u_data_in_ready_prev = '1') then
						cnt <= (cnt + 1);
					end if;
					
					if(cnt < 4) then
						u_valid_in 	<= '1';
						u_data_in 	<= newton_raphson_result((31 - (3-cnt)*8) downto (24 - (3-cnt)*8));
					elsif(cnt < 8) then
						u_valid_in 	<= '1';
						u_data_in 	<= cycle_count((31 - (7-cnt)*8) downto (24 - (7-cnt)*8));
					elsif(cnt < 12) then
						u_valid_in 	<= '1';
						u_data_in 	<= iteration_count((31 - (11-cnt)*8) downto (24 - (11-cnt)*8));
					elsif(cnt < 16) then
						u_valid_in 	<= '1';
						u_data_in 	<= total_cycle_count((31 - (15-cnt)*8) downto (24 - (15-cnt)*8));
					else
						cnt 			<= 0;
						start_opr 	<= '0';
						state			<= power_off;
					end if;
					
				when power_off =>
					leds	 		<= "1000000100";
					state <= reset_all_variable;
					
				when reset_all_variable =>
					state <= idle;
					u_valid_in 					<= '0';
					u_data_in 					<= "01010010";														-- ASCII 'R'
					cnt 							<= 0;
					count							<= 0;
					cycle_count					<= (others => '0');
					total_cycle_count			<= (others => '0');
					degree_min					<= 0;	
					degree_max					<= 0;	
					degree						<= 0;	
					start_opr					<= '0';			
					leds 							<= "0000000000";
					variable_value		  		<= (others => '0');
					float_in(0)  				<= (others => '0');
					float_in(1)  				<= (others => '0');
					float_in(2)  				<= (others => '0');
					float_in(3)  				<= (others => '0');
					float_in(4)  				<= (others => '0');
					float_in(5)  				<= (others => '0');
					float_in(6) 				<= (others => '0');
					float_in(7)  				<= (others => '0');
					float_in(8)  				<= (others => '0');
					float_in(9)  				<= (others => '0');
					float_in(10)  				<= (others => '0');
					float_in(11)				<= (others => '0');
					float_in(12)  				<= (others => '0');
					float_in(13)  				<= (others => '0');
					float_in(14)  				<= (others => '0');
					float_in(15)  				<= (others => '0');
					float_in(16)  				<= (others => '0');
					float_in(17)  				<= (others => '0');
					float_in(18) 				<= (others => '0');
					float_in(19)  				<= (others => '0');
					float_in(20)  				<= (others => '0');
					float_in(21)  				<= (others => '0');
					float_in(22)  				<= (others => '0');
					float_in(23)  				<= (others => '0');
					float_in(24)  				<= (others => '0');
					float_in(25)  				<= (others => '0');
					float_in(26)  				<= (others => '0');
					float_in(27)  				<= (others => '0');
					float_in(28)  				<= (others => '0');
					float_in(29)  				<= (others => '0');
					float_in(30)  				<= (others => '0');
					float_in(31)  				<= (others => '0');
					iteration_count			<= (others => '0');
					error_const_value			<= (others => '0');
					-- End of Program 		
			
				when others =>
					state <= idle;
					
			end case;	
		end if;
	end process;
end logic;	